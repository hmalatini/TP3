`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:29:19 10/31/2016 
// Design Name: 
// Module Name:    Multiplexor_2in_1out 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Multiplexor_2in_1out(
    input [15:0] DatoA,
    input [15:0] DatoB,
    input Sel,
    output reg [15:0] Salida
    );

always @(*)
begin
	if(Sel == 0)
		Salida = DatoA;
	else
		Salida = DatoB;
end

endmodule
